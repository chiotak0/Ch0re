`ifndef CH0RE_TEST_PIPELINE_5ST_SV
`define CH0RE_TEST_PIPELINE_5ST_SV

program tb_pipeline_5st();

endprogram: tb_pipeline_5st

`endif /* CH0RE_TEST_PIPELINE_5ST_SV */
