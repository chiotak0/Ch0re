`include "ch0re_types.sv"





