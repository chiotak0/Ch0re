import ch0re_types::*;

program tb_decoder_id();

    initial begin
        //
    end

endprogram : tb_decoder_id

